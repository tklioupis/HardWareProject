`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:00:25 01/01/2022 
// Design Name: 
// Module Name:    decoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module decoder(
    input [4:0] Awr,
    output [31:0] WEd
    );

	reg [31:0] res;
	assign WEd = res;
	always @(Awr) 
	begin
		case(Awr)
			5'b00000: begin res = 32'b00000000000000000000000000000001; end
			5'b00001: begin res = 32'b00000000000000000000000000000010; end
			5'b00010: begin res = 32'b00000000000000000000000000000100; end
			5'b00011: begin res = 32'b00000000000000000000000000001000; end
			5'b00100: begin res = 32'b00000000000000000000000000010000; end
			5'b00101: begin res = 32'b00000000000000000000000000100000; end
			5'b00110: begin res = 32'b00000000000000000000000001000000; end
			5'b00111: begin res = 32'b00000000000000000000000010000000; end
			5'b01000: begin res = 32'b00000000000000000000000100000000; end			
			5'b01001: begin res = 32'b00000000000000000000001000000000; end
			5'b01010: begin res = 32'b00000000000000000000010000000000; end
			5'b01011: begin res = 32'b00000000000000000000100000000000; end
			5'b01100: begin res = 32'b00000000000000000001000000000000; end
			5'b01101: begin res = 32'b00000000000000000010000000000000; end
			5'b01110: begin res = 32'b00000000000000000100000000000000; end
			5'b01111: begin res = 32'b00000000000000001000000000000000; end
			5'b10000: begin res = 32'b00000000000000010000000000000000; end
			5'b10001: begin res = 32'b00000000000000100000000000000000; end
			5'b10010: begin res = 32'b00000000000001000000000000000000; end
			5'b10011: begin res = 32'b00000000000010000000000000000000; end
			5'b10100: begin res = 32'b00000000000100000000000000000000; end
			5'b10101: begin res = 32'b00000000001000000000000000000000; end
			5'b10110: begin res = 32'b00000000010000000000000000000000; end
			5'b10111: begin res = 32'b00000000100000000000000000000000; end
			5'b11000: begin res = 32'b00000001000000000000000000000000; end
			5'b11001: begin res = 32'b00000010000000000000000000000000; end
			5'b11010: begin res = 32'b00000100000000000000000000000000; end
			5'b11011: begin res = 32'b00001000000000000000000000000000; end
			5'b11100: begin res = 32'b00010000000000000000000000000000; end
			5'b11101: begin res = 32'b00100000000000000000000000000000; end
			5'b11110: begin res = 32'b01000000000000000000000000000000; end
			5'b11111: begin res = 32'b10000000000000000000000000000000; end
		endcase
	end 
endmodule
